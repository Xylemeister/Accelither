
module platform (
	clk_clk,
	filter_in_export,
	reset_reset_n);	

	input		clk_clk;
	input	[15:0]	filter_in_export;
	input		reset_reset_n;
endmodule
